(** * Main module with theorems *)

From ITree Require Export
     Basics.Tacs
     Basics.Basics
     Basics.Category
     Basics.Monad
     Basics.CategoryKleisli
     Basics.CategoryKleisliFacts
     Basics.FunctionFacts
     Core.ITreeDefinition
     Eq
     Core.ITreeMonad
     Core.KTreeFacts
     Indexed.FunctionFacts
     Interp.TranslateFacts
     Interp.InterpFacts
     Interp.HandlerFacts
     Interp.RecursionFacts
     .
